/*******************************************************************
*
* Module: InstMem.v
* Project: Scy_CPU
* Author: Mohamed Sabry momo12320@aucegypt.edu
* Description: Instruction Memory
*
* Change history: 23/10/24 – Reformatted and made to load from a hexfile
*
**********************************************************************/


module InstMem (
 input [9:0] addr,
 output [31:0] data_out
);
reg [31:0] mem [0:(2*1024-1)];
assign data_out = mem[addr];
initial begin
//	mem[0]=32'b0000000000000100000000001_0110111; //LUI
//	mem[1]=32'b0000000000000100000000010_0010111; //AUIPC
//	mem[2]=32'b00000000001000000000000110010011; 
//	mem[3]=32'b00000000010000000000001000010011;
//	mem[4]=32'b11111111111000100000001000010011;
//	mem[5]=32'b00000000010000011000001001100011;
//	mem[6]=32'b00000000000000000000001000010011;
//	mem[7]=32'b00000000001100100001001001100011;
//	mem[8]=32'b00000000000100000000001000010011;
//	mem[9]=32'b00000000001100100001001001100011;
//	mem[10]=32'b00000000011000000000001000010011;
//	mem[11]=32'b00000000001100100100001001100011;
//	mem[12]=32'b00000000011000000000001000010011; //ADDI
//	mem[13]=32'b00000000001100100101001001100011; //BGE
//	mem[14]=32'b00000000001100000000001000010011; //ADDI
//	mem[15]=32'b00000000001100100101001001100011; //BGE
//	mem[16]=32'b00000000001000000000001000010011; //ADDI
//	mem[17]=32'b11111111111000000000001010010011; //ADDI
//	mem[18]=32'b00000000010100100110001001100011; 
//	mem[19]=32'b00000000001000000000001010010011;
//	mem[20]=32'b00000000010000101111001001100011;
//	mem[21]=32'b00000000010000000000001010010011;
//	mem[22]=32'b00000000010000000000001010010011;
//	mem[23]=32'b00000000000000000000000001110011; //ECALL
    /*
    1-addi x1,x0,20	92
    2-addi x2,x0,5	96
    3-add x3,x2,x1	100
    4-jal x5,12(x0)	104
    5-beq x1,x0,126	108
    6-addi x6,x0,1	112
    7-addi x4,x0,0	116
    8-xor x7,x6,x4	120
    9-or x7,x6,x4	124
    10-and x7,x6,x4	128
    11-sub x7,x3,x2	132
    12-slli x7,x2,2	136
    13-slti x7,x2,6	140
    14-addi x8,x0,256565	144
    15-sw x8, 0(x0)	148
    16-sh x8, 4(x0)	152
    17-sb x8, 8(x0)	156
    18-lw x7,0(x0)	160
    19-lh x7,0(x0)	164
    20-lb x7,0(x0)	168
    21-lbu x7,0(x0)	172
    22-lhu x7,0(x0)	176
    23-slti x7,x2,-2	180
    24-xori x7,x2,0	184
    25-ori x7,x2,0	188
    26-andi x7,x2,1	192
    27-srli x7,x2,2	196
    28-srai x7,x2,2	200
    29-addi x9,x0,2	204
    30-sll x7,x2,x9	208
    31-slt x7,x9,x2	212
    32-addi x9,x0,-2	216
    33-sltu x7,x2,x9	220
    34-srl x7,x2,x9	224
    35-sra x7,x2,x9 228
    36-FENCE	232
    37-FENCE.TSO	236
    38-PAUSE	240
    39-addi x1,x0,0	244
    40-JALR x0,0(x5)248
    41-EBREAK	252
    --	
    */
	mem[0]=32'b00000001010000000000000010010011; //addi
	mem[1]=32'b00000000010100000000000100010011; //addi
	mem[2]=32'b00000000000100010000000110110011; //add
	mem[3]=32'b00000000100000000000001011101111; //jal
	mem[4]=32'b00000000000000000000000100010011; //addi
	mem[5]=32'b00000100000000001000100101100011; //beq
	mem[6]=32'b00000000000100000000001100010011; //addi
	mem[7]=32'b00000000000000000000001000010011; // addi
	mem[8]=32'b00000000010000110100001110110011; //xor
	mem[9]=32'b00000000010000110110001110110011; //or
	mem[10]=32'b00000000010000110111001110110011; //and
	mem[11]=32'b01000000001000011000001110110011; //sub
	mem[12]=32'b00000000001000010001001110010011; //slli
	mem[13]=32'b00000000011000010010001110010011; //slti
	
	mem[14]=32'b01111111111100000000010000010011; //addi
	mem[15]=32'b00000000100000000010000000100011; //sw
	mem[16]=32'b00000000100000000001001000100011; //sh
	mem[17]=32'b00000000100000000000010000100011; //sb
	
	mem[18]=32'b00000000000000000100001110000011; //lbu
	mem[19]=32'b00000000000000000000001110000011; //lb
	mem[20]=32'b00000000000000000101001110000011; //lhu
	mem[21]=32'b00000000000000000001001110000011; //lh
    
    
    mem[22]=32'b00000000000000000010001110000011; //lw
	mem[23]=32'b11111111111000010010001110010011; //slti
	mem[24]=32'b00000000000000010100001110010011; //xori
	//         b00000000000000010100001110010011
	mem[25]=32'b00000000000000010110001110010011; //ori
	mem[26]=32'b00000000000100010111001110010011; //andi
	mem[27]=32'b00000000001000010101001110010011; //srli
	mem[28]=32'b01000000001000010101001110010011; //srai
	mem[29]=32'b00000000001000000000010010010011; //addi
	mem[30]=32'b00000000100100010001001110110011; //sll
	mem[31]=32'b00000000001001001010001110110011; //slt
	mem[32]=32'b11111111111000000000010010010011; //addi
	mem[33]=32'b00000000100100010011001110110011; //sltu
	mem[34]=32'b00000000001000000000010010010011; //addi
	
	mem[35]=32'b00000000100100010101001110110011; //srl
	mem[36]=32'b01000000100100010101001110110011; //sra
	mem[37]=32'b0000111111110000000000000_0001111; //fence
	mem[38]=32'b0000000000000000000100000_0001111; //fence.tso
	mem[39]=32'b0000000000000000000100000_0001111; //pause
	mem[40]=32'b00000000000000000000000010010011; //addi 
	mem[41]=32'b00000000000000101000000001100111; //jalr
	mem[42]=32'b00000000000100000000000001110011; //ebreak
	mem[43]=32'b00000000000000000000000001110011; //NOOP
	/*
	00032037
    00032017
    00030313
    00030313
    FFF30313
    00030313
    00030313
    00030313
    00030313
    00030313
    00030313
    00030313
    00030313
    FFF30313
    00030313
    00030313
    00030313
    00030313
	*/
end


endmodule
